module mem(
    
);
    
endmodule