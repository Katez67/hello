module module_1(
    input  a, b, c,
    output sum
);

    assign sum = a + b + c;
    
endmodule