module module_2(
    input  a, b,
    output del
);

    assign del = a - b;
    
endmodule