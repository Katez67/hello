module main(
    input a,
    output b
);

    assign b = a;
    
endmodule